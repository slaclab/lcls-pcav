LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use work.StdRtlPkg.all;

package AppOpts is

  constant APP_TIMING_MODE_C : integer := 1; -- 1 or 2 (LCLS-I/II)
  
end XpmOpts;

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

library surf;
use surf.StdRtlPkg.all;

library xil_default_lib;

package AppOpts is

  constant APP_TIMING_MODE_C : integer := 2; -- 1 or 2 (LCLS-I/II)
  
end AppOpts;
